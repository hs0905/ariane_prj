module reset_ctrl (
  input logic clk,
  input logic rstn,
  input logic state
);
endmodule